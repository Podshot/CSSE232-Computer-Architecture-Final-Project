`timescale 1ns / 1ps

module ProcessorSansControl(
	input clock,
	input MemWrite,
	input [1:0] MemSrc,
	input [2:0] MemDst,
	input [2:0] PCSrc,
	input [1:0] SPSrc,
	input PCWrite,
	input SPWrite,
	input InstWrite,
	input reset,
	input mary_write,
	input shelley_write,
	input comp_write,
	input ra_write,
	input [1:0] mary_src,
	input [1:0] shelley_src,
	input ra_src,
	input SrcA,
	input [1:0] SrcB,
	input [3:0] AluOp,
	input [15:0] io_in,
	output [15:0] io_out,
	output overflow_output,
	output [15:0] instruction
   );

	wire [15:0] mem_out;
	wire [15:0] pc;
	wire [15:0] sp;
	wire [15:0] comp;
	wire [15:0] ra;
	wire [15:0] shelley;
	wire [15:0] mary;
	wire [15:0] sext_imm;
	wire [15:0] sext_ls_imm;
	wire [15:0] zext_imm;
	
	reg [15:0] out_reg;
	reg new_MemWrite;
	reg [15:0] new_MaryData;
	
	always @* begin
		new_MemWrite = MemWrite;
		new_MaryData = mary;
		$display("[PCSP]: MemWrite: %b, MemDst: %b, ze_imm: %b", MemWrite, MemDst, zext_imm);
		if (instruction[14:10] == 5'b10100 && MemWrite == 1 && MemDst == 1 && zext_imm == 255) begin
			out_reg <= mary;
			new_MemWrite = 1'b0;
			$display("[PCSP]: Write to IO -> %b", mary);
			$display("[PCSP]: out_reg: %b", out_reg);
		end
		else if (instruction[14:10] == 5'b10111 && MemWrite == 0 && MemDst == 0 && zext_imm == 255) begin
			$display("[PCSP]: Read from IO");
			new_MaryData = io_in;
		end
		else begin
			out_reg <= 0;
		end
	end
	
	assign io_out = out_reg;

PCSPandMemoryBlock PCSPandMemoryBlock(
	.clock(clock),
	.MemWrite(new_MemWrite),
	.MemSrc(MemSrc),
	.MemDst(MemDst),
	.ze_imm(zext_imm),
	.ls_imm(sext_ls_imm),
	.se_imm(sext_imm),
	.MaryData(mary),
	.ShelleyData(shelley),
	.RAData(ra),
	.CompData(comp),
	.PCSrc(PCSrc),
	.SPSrc(SPSrc),
	.PCWrite(PCWrite),
	.SPWrite(SPWrite),
	.InstWrite(InstWrite),
	.reset(reset),
	.mem_out(mem_out),
	.Inst_out(instruction),
	.pc_out(pc),
	.sp_out(sp)
	);
	
	reg [15:0] inst_reg;
	
	always @ instruction
	begin
		inst_reg = instruction;
	end

RegBlockAndAlu RegBlockAndAlu(
	.memval(mem_out),
	.immediate(inst_reg[9:2]),
	.sp(sp),
	.pc(pc),
	.mary_write(mary_write),
	.shelley_write(shelley_write),
	.comp_write(comp_write),
	.ra_write(ra_write),
	.mary_src(mary_src),
	.shelley_src(shelley_src),
	.ra_src(ra_src),
	.clock(clock),
	.SrcA(SrcA),
	.SrcB(SrcB),
	.AluOp(AluOp),
	.overflow(overflow),
	.mary_output(mary),
	.shelley_output(shelley),
	.comp_output(comp),
	.ra_output(ra),
	.zext_imm_output(zext_imm),
	.sext_imm_output(sext_imm),
	.sext_ls_imm_output(sext_ls_imm),
	.reset(reset)
	);
	
	assign overflow_output = overflow;
	

endmodule
